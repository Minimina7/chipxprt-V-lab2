`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/12/2024 02:17:57 PM
// Design Name: 
// Module Name: tb_addsub4bit
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_addsub4bit;

logic [3:0]a;
logic [3:0]b;
logic cin, Cout; 
logic [3:0] s;
logic M;

addsub4bit result (.a(a), .b(b), .s(s), .CIN(cin), .COUT(Cout), .m(M) );

initial begin

    a[3] = 1'b0;
    a[2] = 1'b0;
    a[1] = 1'b0;
    a[0] = 1'b0;
	b[3] = 1'b0;
	b[2] = 1'b0;
	b[1] = 1'b0;
	b[0] = 1'b0;
	cin = 1'b0;
	M =1'b0;
#5
    a[3] = 1'b0;
    a[2] = 1'b0;
    a[1] = 1'b0;
    a[0] = 1'b1;
	b[3] = 1'b0;
	b[2] = 1'b0;
	b[1] = 1'b0;
	b[0] = 1'b1;
	cin = 1'b0;
	M =1'b1;
#5
    a[3] = 1'b0;
    a[2] = 1'b0;
    a[1] = 1'b1;
    a[0] = 1'b0;
	b[3] = 1'b0;
	b[2] = 1'b0;
	b[1] = 1'b1;
	b[0] = 1'b0;
	cin = 1'b0;
	M =1'b0;
#5
    a[3] = 1'b0;
    a[2] = 1'b0;
    a[1] = 1'b1;
    a[0] = 1'b1;
	b[3] = 1'b0;
	b[2] = 1'b0;
	b[1] = 1'b1;
	b[0] = 1'b1;
	cin = 1'b0;
	M =1'b1;
#5
    a[3] = 1'b0;
    a[2] = 1'b1;
    a[1] = 1'b0;
    a[0] = 1'b0;
	b[3] = 1'b0;
	b[2] = 1'b1;
	b[1] = 1'b0;
	b[0] = 1'b0;
	cin = 1'b0;
	M =1'b0;
#5
    a[3] = 1'b0;
    a[2] = 1'b1;
    a[1] = 1'b0;
    a[0] = 1'b1;
	b[3] = 1'b0;
	b[2] = 1'b1;
	b[1] = 1'b0;
	b[0] = 1'b1;
	cin = 1'b0;
	M =1'b1;
#5
    a[3] = 1'b0;
    a[2] = 1'b1;
    a[1] = 1'b1;
    a[0] = 1'b0;
	b[3] = 1'b0;
	b[2] = 1'b1;
	b[1] = 1'b1;
	b[0] = 1'b0;
	cin = 1'b0;
	M =1'b0;
#5
    a[3] = 1'b0;
    a[2] = 1'b1;
    a[1] = 1'b1;
    a[0] = 1'b1;
	b[3] = 1'b0;
	b[2] = 1'b1;
	b[1] = 1'b1;
	b[0] = 1'b1;
	cin = 1'b0;
	M =1'b1;
#5
    a[3] = 1'b1;
    a[2] = 1'b0;
    a[1] = 1'b0;
    a[0] = 1'b0;
	b[3] = 1'b1;
	b[2] = 1'b0;
	b[1] = 1'b0;
	b[0] = 1'b0;
	cin = 1'b0;
	M =1'b0;
#5
    a[3] = 1'b1;
    a[2] = 1'b0;
    a[1] = 1'b0;
    a[0] = 1'b1;
	b[3] = 1'b1;
	b[2] = 1'b0;
	b[1] = 1'b0;
	b[0] = 1'b1;
	cin = 1'b0;
	M =1'b1;
#5
    a[3] = 1'b1;
    a[2] = 1'b0;
    a[1] = 1'b1;
    a[0] = 1'b0;
	b[3] = 1'b1;
	b[2] = 1'b0;
	b[1] = 1'b1;
	b[0] = 1'b0;
	cin = 1'b0;
	M =1'b0;
#5
    a[3] = 1'b1;
    a[2] = 1'b0;
    a[1] = 1'b1;
    a[0] = 1'b1;
	b[3] = 1'b1;
	b[2] = 1'b0;
	b[1] = 1'b1;
	b[0] = 1'b1;
	cin = 1'b0;
	M =1'b1;
#5
    a[3] = 1'b1;
    a[2] = 1'b1;
    a[1] = 1'b0;
    a[0] = 1'b0;
	b[3] = 1'b1;
	b[2] = 1'b1;
	b[1] = 1'b0;
	b[0] = 1'b0;
	cin = 1'b0;
	M =1'b0;
#5
    a[3] = 1'b1;
    a[2] = 1'b1;
    a[1] = 1'b0;
    a[0] = 1'b1;
	b[3] = 1'b1;
	b[2] = 1'b1;
	b[1] = 1'b0;
	b[0] = 1'b1;
	cin = 1'b0;
	M =1'b1;
#5
    a[3] = 1'b1;
    a[2] = 1'b1;
    a[1] = 1'b1;
    a[0] = 1'b0;
	b[3] = 1'b1;
	b[2] = 1'b1;
	b[1] = 1'b1;
	b[0] = 1'b0;
	cin = 1'b0;
	M =1'b0;
#5
    a[3] = 1'b1;
    a[2] = 1'b1;
    a[1] = 1'b1;
    a[0] = 1'b1;
	b[3] = 1'b1;
	b[2] = 1'b1;
	b[1] = 1'b1;
	b[0] = 1'b1;
	cin = 1'b0;
	M =1'b1;
#5
    a[3] = 1'b0;
    a[2] = 1'b0;
    a[1] = 1'b0;
    a[0] = 1'b0;
	b[3] = 1'b0;
	b[2] = 1'b0;
	b[1] = 1'b0;
	b[0] = 1'b0;
	cin = 1'b1;
	M =1'b0;
#5
    a[3] = 1'b0;
    a[2] = 1'b0;
    a[1] = 1'b0;
    a[0] = 1'b1;
	b[3] = 1'b0;
	b[2] = 1'b0;
	b[1] = 1'b0;
	b[0] = 1'b1;
	cin = 1'b1;
	M =1'b1;
#5
    a[3] = 1'b0;
    a[2] = 1'b0;
    a[1] = 1'b1;
    a[0] = 1'b0;
	b[3] = 1'b0;
	b[2] = 1'b0;
	b[1] = 1'b1;
	b[0] = 1'b0;
	cin = 1'b1;
	M =1'b0;
#5
    a[3] = 1'b0;
    a[2] = 1'b0;
    a[1] = 1'b1;
    a[0] = 1'b1;
	b[3] = 1'b0;
	b[2] = 1'b0;
	b[1] = 1'b1;
	b[0] = 1'b1;
	cin = 1'b1;
	M =1'b1;
#5
    a[3] = 1'b0;
    a[2] = 1'b1;
    a[1] = 1'b0;
    a[0] = 1'b0;
	b[3] = 1'b0;
	b[2] = 1'b1;
	b[1] = 1'b0;
	b[0] = 1'b0;
	cin = 1'b1;
	M =1'b0;
#5
    a[3] = 1'b0;
    a[2] = 1'b1;
    a[1] = 1'b0;
    a[0] = 1'b1;
	b[3] = 1'b0;
	b[2] = 1'b1;
	b[1] = 1'b0;
	b[0] = 1'b1;
	cin = 1'b1;
	M =1'b1;
#5
    a[3] = 1'b0;
    a[2] = 1'b1;
    a[1] = 1'b1;
    a[0] = 1'b0;
	b[3] = 1'b0;
	b[2] = 1'b1;
	b[1] = 1'b1;
	b[0] = 1'b0;
	cin = 1'b1;
	M =1'b0;
#5
    a[3] = 1'b0;
    a[2] = 1'b1;
    a[1] = 1'b1;
    a[0] = 1'b1;
	b[3] = 1'b0;
	b[2] = 1'b1;
	b[1] = 1'b1;
	b[0] = 1'b1;
	cin = 1'b1;
	M =1'b1;
#5
    a[3] = 1'b1;
    a[2] = 1'b0;
    a[1] = 1'b0;
    a[0] = 1'b0;
	b[3] = 1'b1;
	b[2] = 1'b0;
	b[1] = 1'b0;
	b[0] = 1'b0;
	cin = 1'b1;
	M =1'b0;
#5
    a[3] = 1'b1;
    a[2] = 1'b0;
    a[1] = 1'b0;
    a[0] = 1'b1;
	b[3] = 1'b1;
	b[2] = 1'b0;
	b[1] = 1'b0;
	b[0] = 1'b1;
	cin = 1'b1;
	M =1'b1;
#5
    a[3] = 1'b1;
    a[2] = 1'b0;
    a[1] = 1'b1;
    a[0] = 1'b0;
	b[3] = 1'b1;
	b[2] = 1'b0;
	b[1] = 1'b1;
	b[0] = 1'b0;
	cin = 1'b1;
	M =1'b0;
#5
    a[3] = 1'b1;
    a[2] = 1'b0;
    a[1] = 1'b1;
    a[0] = 1'b1;
	b[3] = 1'b1;
	b[2] = 1'b0;
	b[1] = 1'b1;
	b[0] = 1'b1;
	cin = 1'b1;
	M =1'b1;
#5
    a[3] = 1'b1;
    a[2] = 1'b1;
    a[1] = 1'b0;
    a[0] = 1'b0;
	b[3] = 1'b1;
	b[2] = 1'b1;
	b[1] = 1'b0;
	b[0] = 1'b0;
	cin = 1'b1;
	M =1'b0;
#5
    a[3] = 1'b1;
    a[2] = 1'b1;
    a[1] = 1'b0;
    a[0] = 1'b1;
	b[3] = 1'b1;
	b[2] = 1'b1;
	b[1] = 1'b0;
	b[0] = 1'b1;
	cin = 1'b1;
	M =1'b1;
#5
    a[3] = 1'b1;
    a[2] = 1'b1;
    a[1] = 1'b1;
    a[0] = 1'b0;
	b[3] = 1'b1;
	b[2] = 1'b1;
	b[1] = 1'b1;
	b[0] = 1'b0;
	cin = 1'b1;
	M =1'b0;
#5
    a[3] = 1'b1;
    a[2] = 1'b1;
    a[1] = 1'b1;
    a[0] = 1'b1;
	b[3] = 1'b1;
	b[2] = 1'b1;
	b[1] = 1'b1;
	b[0] = 1'b1;
	cin = 1'b1;
	M =1'b1;

#5
$finish;
end

endmodule
